module srt4 (
    input [7:0] inbus,
    input beginSignal, clk, rst_b
    output [7:0] outbus,
    output endSignal
);
    
endmodule